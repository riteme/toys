`ifndef __BPB_VH__
`define __BPB_VH__

`define BPB_E 32
`define BPB_T 11

`endif