`ifndef __CACHE_CONTROLLER_VH__
`define __CACHE_CONTROLLER_VH__

`define NORMAL 4'b1000
`define FETCH 4'b0001
`define WRITE 4'b0000
`define CHECK 4'b0100
`define ALLOC 4'b0010

`endif