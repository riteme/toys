`ifndef __BPB_VH__
`define __BPB_VH__

`define BPB_E 32
`define BPB_T 6

`define T_JMP 0
`define T_JAL 1
`define T_BR 2
`define T_JR 3
`define TMAX `T_JR

// `define USE_BTFNT
// `define USE_GSHARE
// `define USE_LSHARE
`define USE_ALL

`endif