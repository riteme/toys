`ifndef __CACHE_CONTROLLER_VH__
`define __CACHE_CONTROLLER_VH__

`define NORMAL 2'b10
`define FETCH 2'b01
`define WRITE 2'b00

`endif